library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Blink is

    port(    binIn    :    in std_logic_vector(6 downto 0);
            binOut:    out std_logic_vector(6 downto 0);
            clk    :    in std_logic;
            reset    :    in std_logic);

end Blink;

architecture Behavioral of Blink is

    signal last_binIn :    std_logic_vector(6 downto 0);
    signal counter        :    natural;

begin

    process(clk, reset)
    begin
        if(rising_edge(clk)) then    
            if(last_binIn= "1100011" and not (binIn="1100011"))then      
                if(counter=8 or counter=10 or counter=12) then
                    binOut <= (others => '1');
                    counter <= counter+1;
                elsif(counter=7 or counter=9 or counter=11 or counter=13) then
                    binOut <= "1111110";
                    counter <= counter+1;
                else
                    binOut <=(others => '1');
                    counter <= 0;
                end if;
            else
                if(not(last_binIn = binIn)) then
                    last_binIn <= binIn;
                    counter <=0;
                end if;
                
                if(counter=1 or counter=3 or counter=5) then
                    binOut <=(others => '1');
                    counter <= counter+1;
                elsif(counter=0 or counter=2 or counter=4 or counter=6) then
                    binOut <= binIn;
                    counter <= counter+1;
                else
                    binOut <=(others => '1');
                end if;
            end if;
        end if;
    end process;

end Behavioral;