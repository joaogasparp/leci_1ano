library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity SetFSM is
	port(reset : in std_logic;
		  clk : in std_logic;
		  point : in std_logic;
		  seteD : out std_logic;
		  seisD : out std_logic;
		  displayG : out std_logic_vector(6 downto 0));
end SetFSM;

architecture Behav of SetFSM is
	signal s_cntValue : unsigned(2 downto 0);
	type state is (G0, G1, G2, G3, G4, G5, G6, G7);
	signal PS, NS: state;
	constant zeroG : std_logic_vector(6 downto 0) := "1000000"; -- 0
	constant umG : std_logic_vector(6 downto 0) := "1111001"; -- 1
	constant doisG : std_logic_vector(6 downto 0) := "0100100"; -- 2
   constant tresG : std_logic_vector(6 downto 0) := "0110000"; -- 3
   constant quatroG : std_logic_vector(6 downto 0) := "0011001"; -- 4
   constant cincoG : std_logic_vector(6 downto 0) := "0010010"; -- 5
   constant seisG : std_logic_vector(6 downto 0) := "0000010"; -- 6
   constant seteG : std_logic_vector(6 downto 0) := "1111000"; -- 7
begin

   sync_proc : process(clk)
   begin
		if (rising_edge(clk)) then
			if (reset = '0') then
				s_cntValue <= (others => '0');
				PS <= G0;
         elsif (point = '1') then
            s_cntValue <= s_cntValue + 1;
            PS <= NS;
         end if;
		end if;
	end process;

   comb_proc : process(PS, s_cntValue)
   begin
   NS <= PS;

   case PS is
		when G0 =>
			seisD <= '0';
         seteD <= '0';
         displayG <= zeroG;
				
         if (s_cntValue = 1) then
				displayG <= umG;
            NS <= G1;
         end if;

				
		when G1 => 
			if (s_cntValue = 2) then
				displayG <= doisG;
            NS <= G2;
         end if;

			
		when G2 => 
			if (s_cntValue = 3) then
				displayG <= tresG;
            NS <= G3;
         end if;

			
		when G3 =>
			if (s_cntValue = 4) then
				displayG <= quatroG;
            NS <= G4;
         end if;

			
      when G4 =>
         if (s_cntValue = 5) then
				displayG <= cincoG;
            NS <= G5;
         end if;

			
		when G5 =>
			if (s_cntValue = 6) then
				seisD <= '1';
				displayG <= seisG;
            NS <= G6;
			end if;

			
		when G6 =>
			if (s_cntValue = 7) then
				seisD <= '0';
            seteD <= '1';
				displayG <= seteG;
            NS <= G7;
         end if;

			
		when G7 =>
			NS <= G0;
			displayG <= zeroG;

		end case;
	end process;

end Behav;